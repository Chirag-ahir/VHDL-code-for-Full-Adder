-- Testbench for OR gate
library IEEE;
use IEEE.std_logic_1164.all;
 
entity testbench is
-- empty
end testbench; 

architecture tb of testbench is

-- DUT component
component fa1 is
port(
  a: in std_logic;
  b: in std_logic;
  c: in std_logic;
  d: out std_logic;
  e: out std_logic);
end component;


signal a_in, b_in, c_in, d_out,e_out: std_logic;

begin

  -- Connect DUT
  DUT: fa1 port map(a_in, b_in, c_in, d_out,e_out);

  process
  begin
    a_in <= '0';
    b_in <= '0';
    c_in <= '0';
    
    wait for 1 ns;
    
  
     a_in <= '0';
    b_in <= '0';
    c_in <= '1';
  
    wait for 1 ns;
    
    a_in <= '0';
    b_in <= '1';
    c_in <= '0';
    
    wait for 1 ns;
    
    a_in <= '0';
    b_in <= '1';
    c_in <= '1';
    wait for 1 ns;
    
    a_in <= '1';
    b_in <= '0';
    c_in <= '0';
    
    wait for 1 ns;
    
    a_in <= '1';
    b_in <= '0';
    c_in <= '1';
    
    wait for 1 ns;
    
    a_in <= '1';
    b_in <= '1';
    c_in <= '0';
    
    wait for 1 ns;
    
    a_in <= '1';
    b_in <= '1';
    c_in <= '1';
    
    wait for 1 ns;
    
   
    
    wait;
  end process;
end tb;
